App_HW_v0.bsv