// This file is just a catch-all to allow bsc -c to compile all the BC lib files

import  BC_BDPI_decls          :: *;
import  BC_Common              :: *;
import  BC_Dispatch_Adapter    :: *;
import  BC_HW_IFC              :: *;
import  BC_MC_Adapter          :: *;
import  BC_MC_Model            :: *;
import  BC_Management_Adapter  :: *;
import  BC_Mem_Tree            :: *;
import  BC_Transactors         :: *;
import  BC_Utils               :: *;
import  RingNet                :: *;
