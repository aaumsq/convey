App_SSSP.bsv