`ifndef _GALOIS_DEFS_
`define _GALOIS_DEFS_

`define NUM_ENGINES 4
`define NUM_ENGINES_HALF 2
`define LG_NUM_ENGINES 2

//`define WL_SPILL_PORTS 16
//`define WL_WLFIFO_SIZE 1024
`define WL_SPILL_PORTS 16
//`define WL_WLFIFO_SIZE 4

//`define GRAPH_NUM_IN_FLIGHT 192
`define GRAPH_NUM_IN_FLIGHT 256

`define LG_GRAPH_NODE_SIZE 5
`define LG_GRAPH_EDGE_SIZE 3

//`define SSSPENGINE_NUM_IN_FLIGHT 192
//`define SSSPENGINE_NUM_CAS_RETRY_IN_FLIGHT 192
`define SSSPENGINE_NUM_IN_FLIGHT 512
`define SSSPENGINE_NUM_CAS_RETRY_IN_FLIGHT 512

`define WORKLIST_FIFO_SIZE 1024
`define COUNTER_WIDTH 48

`define DEBUG False
`endif
