`ifndef _GALOIS_DEFS_
`define _GALOIS_DEFS_
`define WL_ENGINE_PORTS 16
`define WL_LG_ENGINE_PORTS 4
`define WL_SPILL_PORTS 16
`define WL_WLFIFO_SIZE 1024


`endif