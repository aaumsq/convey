// Copyright (c) 2011-2015 Bluespec, Inc.  All Rights Reserved.
// Distributed under license.

// Author: Rishiyur S. Nikhil

// This package contains some definitions used across the various
// Convey BSV adapters

package BC_Common;

// Some symbolic constants for use in FIFOs to control which interfaces are guarded
Bool ugenq   = True;

Bool ugdeq   = True;

Bool ugcount = True;

endpackage
