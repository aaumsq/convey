`ifndef _GALOIS_DEFS_
`define _GALOIS_DEFS_
`define WL_ENGINE_PORTS 16
`define WL_LG_ENGINE_PORTS 4
`define WL_SPILL_PORTS 16
`define WL_WLFIFO_SIZE 1024

`define GRAPH_PORTS 16
`define GRAPH_NUM_IN_FLIGHT 32

`define LG_GRAPH_NODE_SIZE 4
`define LG_GRAPH_EDGE_SIZE 3

`define DEBUG False
`endif
